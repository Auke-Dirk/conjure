module test_display;
initial begin
  $display ("Let's conjure up a display!");
   #10  $finish;
end
 
endmodule
